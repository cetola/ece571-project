// File: top_hvl.sv
// Authors: 
// Stephano Cetola <cetola@pdx.edu>
//
// Top Level Verification Code
//

`include "definitions.sv"

//use a program block for the testbench
//see 4.3.5 The Program Block and Timing Regions
//Spear, Chris “SystemVerilog for Verification”, Norwell, MA: Springer 2006,
//0-387-27036-1
program top_hvl;

	initial begin

	end

endprogram
